netcdf geopotential_1279l4_0.1x0.1 {
dimensions:
	longitude = 3600 ;
	latitude = 1801 ;
	time = 1 ;
variables:
	float longitude(longitude) ;
		longitude:units = "degrees_east" ;
		longitude:long_name = "longitude" ;
	float latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:long_name = "latitude" ;
	int time(time) ;
		time:units = "hours since 1900-01-01 00:00:00.0" ;
		time:long_name = "time" ;
		time:calendar = "gregorian" ;
	short z(time, latitude, longitude) ;
		z:scale_factor = 1.00450154883799 ;
		z:add_offset = 29342.9235304756 ;
		z:_FillValue = -32767s ;
		z:missing_value = -32767s ;
		z:units = "m**2 s**-2" ;
		z:long_name = "Geopotential" ;
		z:standard_name = "geopotential" ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:history = "2020-05-28 21:39:20 GMT by grib_to_netcdf-2.16.0: grib_to_netcdf -o geopotential_1279l4_0.1x0.1.nc geo_1279l4_0.1x0.1.grb" ;
}
